----------------------------------------------------------------------------------
--Ben Oztalay, 2009-2010
--
--This VHDL code is part of the OZ-3, a 32-bit processor
--
--Module Title: EX
--Module Description:
--	The Execution stage of the OZ-3, which performs all of the arithmetic,
-- generates the flags for use with branch instructions, and ultimately makes
-- the choice to branch or not.
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity EX is
	Port ( clock : in STD_LOGIC;
		    reset : in STD_LOGIC;
			 ALUA_from_ID  : in STD_LOGIC_VECTOR(31 downto 0);
			 ALUB_from_ID  : in STD_LOGIC_VECTOR(31 downto 0);
			 cntl_from_ID : in STD_LOGIC_VECTOR(11 downto 0);
			 p_flag_from_MEM : in STD_LOGIC;
			 ALUR_to_MEM : out STD_LOGIC_VECTOR(31 downto 0);
			 dest_reg_addr_to_ID : out STD_LOGIC_VECTOR(4 downto 0);
			 cond_bit_to_IF : out STD_LOGIC);
end EX;

architecture Behavioral of EX is

--//Components\\--

--The Arithmetic and Logic Unit
component ALU is
    Port ( A : in  STD_LOGIC_VECTOR (31 downto 0);
           B : in  STD_LOGIC_VECTOR (31 downto 0);
           sel : in  STD_LOGIC_VECTOR (3 downto 0);
           result : out  STD_LOGIC_VECTOR (31 downto 0);
           flags : out  STD_LOGIC_VECTOR (3 downto 0));
end component;

--The condition block, which holds all of the flags generated by the
--ALU and sends the selected flag to the IF stage
component ConditionBlock is
	Port ( clock : in STD_LOGIC;
			 reset : in STD_LOGIC;
			 sel   : in STD_LOGIC_VECTOR(2 downto 0);
			 flags : in STD_LOGIC_VECTOR(4 downto 0);
			 cond_out : out STD_LOGIC);
end component;

--Generic rising-edge-triggered register
component GenReg is
	 generic (size: integer);
		 Port ( clock : in  STD_LOGIC;
				  enable : in STD_LOGIC;
				  reset : in  STD_LOGIC;
				  data : in  STD_LOGIC_VECTOR ((size - 1) downto 0);
				  output : out  STD_LOGIC_VECTOR ((size - 1) downto 0));
end component;

--\\Components//--

--//Signals\\--

signal ALUA_reg_out : STD_LOGIC_VECTOR(31 downto 0); --Output of the stage's input registers
signal ALUB_reg_out : STD_LOGIC_VECTOR(31 downto 0); 
signal ALU_flags    : STD_LOGIC_VECTOR(3 downto 0);  --Carries the flags generated by the ALU
signal cntl_reg_out : STD_LOGIC_VECTOR(11 downto 0); --This is the output of the 1-stage buffer that delays the
																	  --control signals coming from the decoder
signal flags_to_CB  : STD_LOGIC_VECTOR(4 downto 0);  --Carries all of the flags to the condition block, including
																	  --the pin flag from MEMIO
--\\Signals//--

begin

	--ALU instantiation
	ALU_inst: ALU port map (A => ALUA_reg_out,
									B => ALUB_reg_out,
									sel => cntl_reg_out(3 downto 0),
									result => ALUR_to_MEM,
									flags => ALU_flags);
	
	--Condition Block instantiation
	cond_block: ConditionBlock port map (clock => clock, 
													 reset => reset, 
													 sel => cntl_reg_out(6 downto 4),
													 flags => flags_to_CB,
													 cond_out => cond_bit_to_IF);

	--Input register A instantiation
	ALUA_reg: GenReg generic map (size => 32)
	                 port map (clock => clock,
										enable => '1',
										reset => reset,
										data => ALUA_from_ID,
										output => ALUA_reg_out);
										
	--Input register B instantiation
	ALUB_reg: GenReg generic map (size => 32)
	                 port map (clock => clock,
										enable => '1', 
										reset => reset, 
										data => ALUB_from_ID, 
										output => ALUB_reg_out);
										
	--Control signal buffer register 1 instantiation
	Cntl_reg: GenReg generic map (size => 12)
						  port map (clock => clock, 
										enable => '1', 
										reset => reset, 
										data => cntl_from_ID, 
										output => cntl_reg_out);
						  
	flags_to_CB <= (p_flag_from_MEM & ALU_flags); --Adding the pin flag to the ALU flags
	dest_reg_addr_to_ID <= cntl_reg_out(11 downto 7); --Sending the instruction's result register back to ID for
end Behavioral;												  --forwarding logic

